module icache(
    
    );
endmodule
